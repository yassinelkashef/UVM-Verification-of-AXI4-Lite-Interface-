package AXI_pkg;


 import uvm_pkg::*;
 
 `include "uvm_macros.svh"
  



  `include "Seq_Item.sv"
  `include "Sequencer.sv"
  `include "Monitor.sv"
  `include "Driver.sv"
  `include "Coverage_Collector.sv"
  `include "Agent.sv"
  `include "Environment.sv"
  `include "Base_Sequence.sv"
  `include "AXI_Reset_Seq.sv"
  `include "AXI_Write_Data_8.sv"
  `include "AXI_Write_Data_16.sv"
  `include "AXI_Write_Data_32.sv"
  `include "AXI_Read_Data.sv"
  `include "AXI_Test.sv"
 



endpackage 
